//----------------------------------------------------------------------------------------------------
// Filename: IF_Stage_tb.sv
// Author: Charles Bassani
// Description: Testbench for IF_Stage
//----------------------------------------------------------------------------------------------------
`timescale 1ns/1ps

//----------------------------------------------------------------------------------------------------
// Module Declaration
//----------------------------------------------------------------------------------------------------
module IF_Stage_tb;

//----------------------------------------------------------------------------------------------------
// Test Registers
//----------------------------------------------------------------------------------------------------
logic        clk;
logic        rst;
logic        stall;
logic        flush;
logic [31:0] pc_in;
logic [31:0] pc_out;
logic [31:0] instruction_out;

//----------------------------------------------------------------------------------------------------
// Device Under Test
//----------------------------------------------------------------------------------------------------
IF_Stage dut
(
    .clk(clk),
    .rst(rst),
    .stall(stall),
    .flush(flush),
    .pc_in(pc_in),
    .pc_out(pc_out),
    .instruction_out(instruction_out)
);

//----------------------------------------------------------------------------------------------------
// Waveform Generation
//----------------------------------------------------------------------------------------------------
initial begin
    $dumpfile("build/IF_Stage_tb_wave.vcd");
    $dumpvars(0, IF_Stage_tb);
end

//----------------------------------------------------------------------------------------------------
// Memory Load
//----------------------------------------------------------------------------------------------------
initial begin
    string filename;
    if(!$value$plusargs("IMEM_FILE=%s", filename)) filename = "programs/imem_init.hex";
    $readmemh(filename, dut.imem_inst.mem);
end

//----------------------------------------------------------------------------------------------------
// Test Logic
//----------------------------------------------------------------------------------------------------
always #5 clk = ~clk;

initial begin
    //Initialize signals
    clk   = 0;
    rst   = 1;
    stall = 0;
    flush = 0;
    pc_in = 32'b0;

    //Hold reset for a few cycles
    #10 rst = 0;

    //Increment PC
    for(int i = 0; i < 25; ++i) begin
        pc_in = pc_in + 4; 
        #10 $display("PC: %x, Instruction: %x", pc_out, instruction_out);
    end

    $finish;
end

endmodule
